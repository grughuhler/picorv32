/* Copyright 2024 Grug Huhler.  License SPDX BSD-2-Clause. */

// 8192 bytes of sram formed from 4 Gowin single-port BSRAMs.

module sram
  #(parameter ADDRWIDTH=13)
   (
    input wire                 clk,
    input wire                 resetn,
    input wire                 sram_sel,
    input wire [3:0]           wstrb,
    input wire [ADDRWIDTH-1:0] addr,
    input wire [31:0]          sram_data_i,
    output wire                sram_ready,
    output wire [31:0]         sram_data_o
    );
 
   // This is the memory initialization file formed by program conv_to_init.
   // Be sure this file rebuilds if the include file is changed.
   `include "mem_init.v"

   reg ready = 1'b0;

   assign sram_ready = ready;
   
   Gowin_SP #(
              .INIT_RAM_00(RAM3_00),
              .INIT_RAM_01(RAM3_01),
              .INIT_RAM_02(RAM3_02),
              .INIT_RAM_03(RAM3_03),
              .INIT_RAM_04(RAM3_04),
              .INIT_RAM_05(RAM3_05),
              .INIT_RAM_06(RAM3_06),
              .INIT_RAM_07(RAM3_07),
              .INIT_RAM_08(RAM3_08),
              .INIT_RAM_09(RAM3_09),
              .INIT_RAM_0A(RAM3_0A),
              .INIT_RAM_0B(RAM3_0B),
              .INIT_RAM_0C(RAM3_0C),
              .INIT_RAM_0D(RAM3_0D),
              .INIT_RAM_0E(RAM3_0E),
              .INIT_RAM_0F(RAM3_0F),
              .INIT_RAM_10(RAM3_10),
              .INIT_RAM_11(RAM3_11),
              .INIT_RAM_12(RAM3_12),
              .INIT_RAM_13(RAM3_13),
              .INIT_RAM_14(RAM3_14),
              .INIT_RAM_15(RAM3_15),
              .INIT_RAM_16(RAM3_16),
              .INIT_RAM_17(RAM3_17),
              .INIT_RAM_18(RAM3_18),
              .INIT_RAM_19(RAM3_19),
              .INIT_RAM_1A(RAM3_1A),
              .INIT_RAM_1B(RAM3_1B),
              .INIT_RAM_1C(RAM3_1C),
              .INIT_RAM_1D(RAM3_1D),
              .INIT_RAM_1E(RAM3_1E),
              .INIT_RAM_1F(RAM3_1F),
              .INIT_RAM_20(RAM3_20),
              .INIT_RAM_21(RAM3_21),
              .INIT_RAM_22(RAM3_22),
              .INIT_RAM_23(RAM3_23),
              .INIT_RAM_24(RAM3_24),
              .INIT_RAM_25(RAM3_25),
              .INIT_RAM_26(RAM3_26),
              .INIT_RAM_27(RAM3_27),
              .INIT_RAM_28(RAM3_28),
              .INIT_RAM_29(RAM3_29),
              .INIT_RAM_2A(RAM3_2A),
              .INIT_RAM_2B(RAM3_2B),
              .INIT_RAM_2C(RAM3_2C),
              .INIT_RAM_2D(RAM3_2D),
              .INIT_RAM_2E(RAM3_2E),
              .INIT_RAM_2F(RAM3_2F),
              .INIT_RAM_30(RAM3_30),
              .INIT_RAM_31(RAM3_31),
              .INIT_RAM_32(RAM3_32),
              .INIT_RAM_33(RAM3_33),
              .INIT_RAM_34(RAM3_34),
              .INIT_RAM_35(RAM3_35),
              .INIT_RAM_36(RAM3_36),
              .INIT_RAM_37(RAM3_37),
              .INIT_RAM_38(RAM3_38),
              .INIT_RAM_39(RAM3_39),
              .INIT_RAM_3A(RAM3_3A),
              .INIT_RAM_3B(RAM3_3B),
              .INIT_RAM_3C(RAM3_3C),
              .INIT_RAM_3D(RAM3_3D),
              .INIT_RAM_3E(RAM3_3E),
              .INIT_RAM_3F(RAM3_3F)
              )
   gmem3
     (
      .dout(sram_data_o[31:24]),
      .clk(clk),
      .oce(1'b1),
      .ce(sram_sel),
      .reset(~resetn),
      .wre(wstrb[3]),
      .ad(addr[12:2]),
      .din(sram_data_i[31:24])
      );

   Gowin_SP #(
              .INIT_RAM_00(RAM2_00),
              .INIT_RAM_01(RAM2_01),
              .INIT_RAM_02(RAM2_02),
              .INIT_RAM_03(RAM2_03),
              .INIT_RAM_04(RAM2_04),
              .INIT_RAM_05(RAM2_05),
              .INIT_RAM_06(RAM2_06),
              .INIT_RAM_07(RAM2_07),
              .INIT_RAM_08(RAM2_08),
              .INIT_RAM_09(RAM2_09),
              .INIT_RAM_0A(RAM2_0A),
              .INIT_RAM_0B(RAM2_0B),
              .INIT_RAM_0C(RAM2_0C),
              .INIT_RAM_0D(RAM2_0D),
              .INIT_RAM_0E(RAM2_0E),
              .INIT_RAM_0F(RAM2_0F),
              .INIT_RAM_10(RAM2_10),
              .INIT_RAM_11(RAM2_11),
              .INIT_RAM_12(RAM2_12),
              .INIT_RAM_13(RAM2_13),
              .INIT_RAM_14(RAM2_14),
              .INIT_RAM_15(RAM2_15),
              .INIT_RAM_16(RAM2_16),
              .INIT_RAM_17(RAM2_17),
              .INIT_RAM_18(RAM2_18),
              .INIT_RAM_19(RAM2_19),
              .INIT_RAM_1A(RAM2_1A),
              .INIT_RAM_1B(RAM2_1B),
              .INIT_RAM_1C(RAM2_1C),
              .INIT_RAM_1D(RAM2_1D),
              .INIT_RAM_1E(RAM2_1E),
              .INIT_RAM_1F(RAM2_1F),
              .INIT_RAM_20(RAM2_20),
              .INIT_RAM_21(RAM2_21),
              .INIT_RAM_22(RAM2_22),
              .INIT_RAM_23(RAM2_23),
              .INIT_RAM_24(RAM2_24),
              .INIT_RAM_25(RAM2_25),
              .INIT_RAM_26(RAM2_26),
              .INIT_RAM_27(RAM2_27),
              .INIT_RAM_28(RAM2_28),
              .INIT_RAM_29(RAM2_29),
              .INIT_RAM_2A(RAM2_2A),
              .INIT_RAM_2B(RAM2_2B),
              .INIT_RAM_2C(RAM2_2C),
              .INIT_RAM_2D(RAM2_2D),
              .INIT_RAM_2E(RAM2_2E),
              .INIT_RAM_2F(RAM2_2F),
              .INIT_RAM_30(RAM2_30),
              .INIT_RAM_31(RAM2_31),
              .INIT_RAM_32(RAM2_32),
              .INIT_RAM_33(RAM2_33),
              .INIT_RAM_34(RAM2_34),
              .INIT_RAM_35(RAM2_35),
              .INIT_RAM_36(RAM2_36),
              .INIT_RAM_37(RAM2_37),
              .INIT_RAM_38(RAM2_38),
              .INIT_RAM_39(RAM2_39),
              .INIT_RAM_3A(RAM2_3A),
              .INIT_RAM_3B(RAM2_3B),
              .INIT_RAM_3C(RAM2_3C),
              .INIT_RAM_3D(RAM2_3D),
              .INIT_RAM_3E(RAM2_3E),
              .INIT_RAM_3F(RAM2_3F)
              )
     gmem2
     (
      .dout(sram_data_o[23:16]),
      .clk(clk),
      .oce(1'b1),
      .ce(sram_sel),
      .reset(~resetn),
      .wre(wstrb[2]),
      .ad(addr[12:2]),
      .din(sram_data_i[23:16])
      );

   Gowin_SP #(
              .INIT_RAM_00(RAM1_00),
              .INIT_RAM_01(RAM1_01),
              .INIT_RAM_02(RAM1_02),
              .INIT_RAM_03(RAM1_03),
              .INIT_RAM_04(RAM1_04),
              .INIT_RAM_05(RAM1_05),
              .INIT_RAM_06(RAM1_06),
              .INIT_RAM_07(RAM1_07),
              .INIT_RAM_08(RAM1_08),
              .INIT_RAM_09(RAM1_09),
              .INIT_RAM_0A(RAM1_0A),
              .INIT_RAM_0B(RAM1_0B),
              .INIT_RAM_0C(RAM1_0C),
              .INIT_RAM_0D(RAM1_0D),
              .INIT_RAM_0E(RAM1_0E),
              .INIT_RAM_0F(RAM1_0F),
              .INIT_RAM_10(RAM1_10),
              .INIT_RAM_11(RAM1_11),
              .INIT_RAM_12(RAM1_12),
              .INIT_RAM_13(RAM1_13),
              .INIT_RAM_14(RAM1_14),
              .INIT_RAM_15(RAM1_15),
              .INIT_RAM_16(RAM1_16),
              .INIT_RAM_17(RAM1_17),
              .INIT_RAM_18(RAM1_18),
              .INIT_RAM_19(RAM1_19),
              .INIT_RAM_1A(RAM1_1A),
              .INIT_RAM_1B(RAM1_1B),
              .INIT_RAM_1C(RAM1_1C),
              .INIT_RAM_1D(RAM1_1D),
              .INIT_RAM_1E(RAM1_1E),
              .INIT_RAM_1F(RAM1_1F),
              .INIT_RAM_20(RAM1_20),
              .INIT_RAM_21(RAM1_21),
              .INIT_RAM_22(RAM1_22),
              .INIT_RAM_23(RAM1_23),
              .INIT_RAM_24(RAM1_24),
              .INIT_RAM_25(RAM1_25),
              .INIT_RAM_26(RAM1_26),
              .INIT_RAM_27(RAM1_27),
              .INIT_RAM_28(RAM1_28),
              .INIT_RAM_29(RAM1_29),
              .INIT_RAM_2A(RAM1_2A),
              .INIT_RAM_2B(RAM1_2B),
              .INIT_RAM_2C(RAM1_2C),
              .INIT_RAM_2D(RAM1_2D),
              .INIT_RAM_2E(RAM1_2E),
              .INIT_RAM_2F(RAM1_2F),
              .INIT_RAM_30(RAM1_30),
              .INIT_RAM_31(RAM1_31),
              .INIT_RAM_32(RAM1_32),
              .INIT_RAM_33(RAM1_33),
              .INIT_RAM_34(RAM1_34),
              .INIT_RAM_35(RAM1_35),
              .INIT_RAM_36(RAM1_36),
              .INIT_RAM_37(RAM1_37),
              .INIT_RAM_38(RAM1_38),
              .INIT_RAM_39(RAM1_39),
              .INIT_RAM_3A(RAM1_3A),
              .INIT_RAM_3B(RAM1_3B),
              .INIT_RAM_3C(RAM1_3C),
              .INIT_RAM_3D(RAM1_3D),
              .INIT_RAM_3E(RAM1_3E),
              .INIT_RAM_3F(RAM1_3F)
              )
     gmem1
     (
      .dout(sram_data_o[15:8]),
      .clk(clk),
      .oce(1'b1),
      .ce(sram_sel),
      .reset(~resetn),
      .wre(wstrb[1]),
      .ad(addr[12:2]),
      .din(sram_data_i[15:8])
      );

   Gowin_SP #(
              .INIT_RAM_00(RAM0_00),
              .INIT_RAM_01(RAM0_01),
              .INIT_RAM_02(RAM0_02),
              .INIT_RAM_03(RAM0_03),
              .INIT_RAM_04(RAM0_04),
              .INIT_RAM_05(RAM0_05),
              .INIT_RAM_06(RAM0_06),
              .INIT_RAM_07(RAM0_07),
              .INIT_RAM_08(RAM0_08),
              .INIT_RAM_09(RAM0_09),
              .INIT_RAM_0A(RAM0_0A),
              .INIT_RAM_0B(RAM0_0B),
              .INIT_RAM_0C(RAM0_0C),
              .INIT_RAM_0D(RAM0_0D),
              .INIT_RAM_0E(RAM0_0E),
              .INIT_RAM_0F(RAM0_0F),
              .INIT_RAM_10(RAM0_10),
              .INIT_RAM_11(RAM0_11),
              .INIT_RAM_12(RAM0_12),
              .INIT_RAM_13(RAM0_13),
              .INIT_RAM_14(RAM0_14),
              .INIT_RAM_15(RAM0_15),
              .INIT_RAM_16(RAM0_16),
              .INIT_RAM_17(RAM0_17),
              .INIT_RAM_18(RAM0_18),
              .INIT_RAM_19(RAM0_19),
              .INIT_RAM_1A(RAM0_1A),
              .INIT_RAM_1B(RAM0_1B),
              .INIT_RAM_1C(RAM0_1C),
              .INIT_RAM_1D(RAM0_1D),
              .INIT_RAM_1E(RAM0_1E),
              .INIT_RAM_1F(RAM0_1F),
              .INIT_RAM_20(RAM0_20),
              .INIT_RAM_21(RAM0_21),
              .INIT_RAM_22(RAM0_22),
              .INIT_RAM_23(RAM0_23),
              .INIT_RAM_24(RAM0_24),
              .INIT_RAM_25(RAM0_25),
              .INIT_RAM_26(RAM0_26),
              .INIT_RAM_27(RAM0_27),
              .INIT_RAM_28(RAM0_28),
              .INIT_RAM_29(RAM0_29),
              .INIT_RAM_2A(RAM0_2A),
              .INIT_RAM_2B(RAM0_2B),
              .INIT_RAM_2C(RAM0_2C),
              .INIT_RAM_2D(RAM0_2D),
              .INIT_RAM_2E(RAM0_2E),
              .INIT_RAM_2F(RAM0_2F),
              .INIT_RAM_30(RAM0_30),
              .INIT_RAM_31(RAM0_31),
              .INIT_RAM_32(RAM0_32),
              .INIT_RAM_33(RAM0_33),
              .INIT_RAM_34(RAM0_34),
              .INIT_RAM_35(RAM0_35),
              .INIT_RAM_36(RAM0_36),
              .INIT_RAM_37(RAM0_37),
              .INIT_RAM_38(RAM0_38),
              .INIT_RAM_39(RAM0_39),
              .INIT_RAM_3A(RAM0_3A),
              .INIT_RAM_3B(RAM0_3B),
              .INIT_RAM_3C(RAM0_3C),
              .INIT_RAM_3D(RAM0_3D),
              .INIT_RAM_3E(RAM0_3E),
              .INIT_RAM_3F(RAM0_3F)
              )
     gmem0
     (
      .dout(sram_data_o[7:0]),
      .clk(clk),
      .oce(1'b1),
      .ce(sram_sel),
      .reset(~resetn),
      .wre(wstrb[0]),
      .ad(addr[12:2]),
      .din(sram_data_i[7:0])
      );

   always @(posedge clk) 
     if (sram_sel)
        ready <= 1'b1;
     else
        ready <= 1'b0;


   
endmodule // sram
